// ==================================================
// Copyright (c)
// All rights reserved
// Filename        : riscv_dut.sv
// Author          : x00897025
// Email           : 1834093202@qq.com
// Created on      : 2024-11-23 03:38:22
// Last Modified   : 2024-11-23 04:30:01
// Description     : 
// 
// 
// ==================================================

